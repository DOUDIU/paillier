/*
    X = x10x9x8x7x6x5x4x3x2x1x0
    Y = y7y6y5y4y3y2yy15y14y13y12y11y10y9y8y7y6y5y4y3y2y1y01y0
    X*Y = (x10x9x8x7x6x5x4x3x2x1x0) * (y15y14y13y12y11y10y9y8y7y6y5y4y3y2y1y0)
        = ((x10 << 240) + (x9 << 216) + (x8 << 192) + (x7 << 168) + (x6 << 144) + (x5 << 120) + (x4 << 96) + (x3 << 72) + (x2 << 48) + (x1 << 24) + x0)
            * ((y15 << 240) + (y14 << 224) + (y13 << 208) + (y12 << 192) + (y11 << 176) + (y10 << 160) + (y9 << 144) + (y8 << 128) + (y7 << 112) + (y6 << 96) + (y5 << 80) + (y4 << 64) + (y3 << 48) + (y2 << 32) + (y1 << 16) + y0)
        =  (
            (x10y15) << 480
        +   (x10y14) << 464
        +   (x9y15 ) << 456
        +   (x10y13) << 448
        +   (x9y14 ) << 440
        +   (x10y12) << 432
        +   (x8y15 ) << 432
        +   (x9y13 ) << 424
        +   (x10y11) << 416
        +   (x8y14 ) << 416
        +   (x9y12 ) << 408
        +   (x7y15 ) << 408
        +   (x10y10) << 400
        +   (x8y13 ) << 400
        +   (x9y11 ) << 392
        +   (x7y14 ) << 392
        +   (x10y9 ) << 384
        +   (x8y12 ) << 384
        +   (x6y15 ) << 384
        +   (x9y10 ) << 376
        +   (x7y13 ) << 376
        +   (x10y8 ) << 368
        +   (x8y11 ) << 368
        +   (x6y14 ) << 368
        +   (x9y9  ) << 360
        +   (x7y12 ) << 360
        +   (x5y15 ) << 360
        +   (x10y7 ) << 352
        +   (x8y10 ) << 352
        +   (x6y13 ) << 352
        +   (x9y8  ) << 344
        +   (x7y11 ) << 344
        +   (x5y14 ) << 344
        +   (x10y6 ) << 336
        +   (x8y9  ) << 336
        +   (x6y12 ) << 336
        +   (x4y15 ) << 336
        +   (x9y7  ) << 328
        +   (x7y10 ) << 328
        +   (x5y13 ) << 328
        +   (x10y5 ) << 320
        +   (x8y8  ) << 320
        +   (x6y11 ) << 320
        +   (x4y14 ) << 320
        +   (x9y6  ) << 312
        +   (x7y9  ) << 312
        +   (x5y12 ) << 312
        +   (x3y15 ) << 312
        +   (x10y4 ) << 304
        +   (x8y7  ) << 304
        +   (x6y10 ) << 304
        +   (x4y13 ) << 304
        +   (x9y5  ) << 296
        +   (x7y8  ) << 296
        +   (x5y11 ) << 296
        +   (x3y14 ) << 296
        +   (x10y3 ) << 288
        +   (x8y6  ) << 288
        +   (x6y9  ) << 288
        +   (x4y12 ) << 288
        +   (x2y15 ) << 288
        +   (x9y4  ) << 280
        +   (x7y7  ) << 280
        +   (x5y10 ) << 280
        +   (x3y13 ) << 280
        +   (x10y2 ) << 272
        +   (x8y5  ) << 272
        +   (x6y8  ) << 272
        +   (x4y11 ) << 272
        +   (x2y14 ) << 272
        +   (x9y3  ) << 264
        +   (x7y6  ) << 264
        +   (x5y9  ) << 264
        +   (x3y12 ) << 264
        +   (x1y15 ) << 264
        +   (x10y1 ) << 256
        +   (x8y4  ) << 256
        +   (x6y7  ) << 256
        +   (x4y10 ) << 256
        +   (x2y13 ) << 256
        +   (x9y2  ) << 248
        +   (x7y5  ) << 248
        +   (x5y8  ) << 248
        +   (x3y11 ) << 248
        +   (x1y14 ) << 248
        +   (x10y0 ) << 240
        +   (x8y3  ) << 240
        +   (x6y6  ) << 240
        +   (x4y9  ) << 240
        +   (x2y12 ) << 240
        +   (x0y15 ) << 240
        +   (x9y1  ) << 232
        +   (x7y4  ) << 232
        +   (x5y7  ) << 232
        +   (x3y10 ) << 232
        +   (x1y13 ) << 232
        +   (x8y2  ) << 224
        +   (x6y5  ) << 224
        +   (x4y8  ) << 224
        +   (x0y14 ) << 224
        +   (x2y11 ) << 224
        +   (x9y0  ) << 216
        +   (x7y3  ) << 216
        +   (x5y6  ) << 216
        +   (x3y9  ) << 216
        +   (x1y12 ) << 216
        +   (x8y1  ) << 208
        +   (x6y4  ) << 208
        +   (x4y7  ) << 208
        +   (x2y10 ) << 208
        +   (x0y13 ) << 208
        +   (x7y2  ) << 200
        +   (x5y5  ) << 200
        +   (x3y8  ) << 200
        +   (x1y11 ) << 200
        +   (x8y0  ) << 192
        +   (x6y3  ) << 192
        +   (x4y6  ) << 192
        +   (x2y9  ) << 192
        +   (x0y12 ) << 192
        +   (x7y1  ) << 184
        +   (x5y4  ) << 184
        +   (x3y7  ) << 184
        +   (x1y10 ) << 184
        +   (x6y2  ) << 176
        +   (x4y5  ) << 176
        +   (x2y8  ) << 176
        +   (x0y11 ) << 176
        +   (x7y0  ) << 168
        +   (x5y3  ) << 168
        +   (x3y6  ) << 168
        +   (x1y9  ) << 168
        +   (x6y1  ) << 160
        +   (x4y4  ) << 160
        +   (x2y7  ) << 160
        +   (x0y10 ) << 160
        +   (x5y2  ) << 152
        +   (x3y5  ) << 152
        +   (x1y8  ) << 152
        +   (x6y0  ) << 144
        +   (x4y3  ) << 144
        +   (x2y6  ) << 144
        +   (x0y9  ) << 144
        +   (x5y1  ) << 136
        +   (x3y4  ) << 136
        +   (x1y7  ) << 136
        +   (x4y2  ) << 128
        +   (x2y5  ) << 128
        +   (x0y8  ) << 128
        +   (x5y0  ) << 120
        +   (x3y3  ) << 120
        +   (x1y6  ) << 120
        +   (x4y1  ) << 112
        +   (x2y4  ) << 112
        +   (x0y7  ) << 112
        +   (x3y2  ) << 104
        +   (x1y5  ) << 104
        +   (x4y0  ) << 96
        +   (x2y3  ) << 96
        +   (x0y6  ) << 96
        +   (x3y1  ) << 88
        +   (x1y4  ) << 88
        +   (x0y5  ) << 80
        +   (x2y2  ) << 80
        +   (x3y0  ) << 72
        +   (x1y3  ) << 72
        +   (x2y1  ) << 64
        +   (x0y4  ) << 64
        +   (x1y2  ) << 56
        +   (x2y0  ) << 48
        +   (x0y3  ) << 48
        +   (x1y1  ) << 40
        +   (x0y2  ) << 32
        +   (x1y0  ) << 24
        +   (x0y1  ) << 16
        +   (x0y0  )
    )
*/
/*
    X = x10x9x8x7x6x5x4x3x2x1x0
    Y = y7y6y5y4y3y2yy15y14y13y12y11y10y9y8y7y6y5y4y3y2y1y01y0
    X*Y = (x10x9x8x7x6x5x4x3x2x1x0) * (y15y14y13y12y11y10y9y8y7y6y5y4y3y2y1y0)
        = ((x10 << 240) + (x9 << 216) + (x8 << 192) + (x7 << 168) + (x6 << 144) + (x5 << 120) + (x4 << 96) + (x3 << 72) + (x2 << 48) + (x1 << 24) + x0)
            * ((y15 << 240) + (y14 << 224) + (y13 << 208) + (y12 << 192) + (y11 << 176) + (y10 << 160) + (y9 << 144) + (y8 << 128) + (y7 << 112) + (y6 << 96) + (y5 << 80) + (y4 << 64) + (y3 << 48) + (y2 << 32) + (y1 << 16) + y0)
        =  (
            (x10y15) << 480
        +   (x10y14) << 464
        +   (x9y15 ) << 456
        +   (x10y13) << 448
        +   (x9y14 ) << 440
        +   (x8y15 + x10y12) << 432
        +   (x9y13 ) << 424
        +   (x8y14 + x10y11) << 416
        +   (x7y15 + x9y12) << 408
        +   (x8y13 + x10y10) << 400
        +   (x7y14 + x9y11) << 392
        +   (x6y15 + x8y12 + x10y9) << 384

        +   (x7y13 + x9y10) << 376
        +   (x6y14 + x8y11 + x10y8) << 368
        +   (x5y15 + x7y12 + x9y9) << 360
        +   (x6y13 + x8y10 + x10y7) << 352
        +   (x5y14 + x7y11 + x9y8) << 344
        +   (x4y15 + x6y12 + x8y9 + x10y6) << 336
        +   (x5y13 + x7y10 + x9y7) << 328
        +   (x4y14 + x6y11 + x8y8 + x10y5) << 320
        +   (x3y15 + x5y12 + x7y9 + x9y6) << 312
        +   (x4y13 + x6y10 + x8y7 + x10y4) << 304
        +   (x3y14 + x5y11 + x7y8 + x9y5) << 296
        +   (x2y15 + x4y12 + x6y9 + x8y6 + x10y3) << 288
        +   (x3y13 + x5y10 + x7y7 + x9y4) << 280
        +   (x2y14 + x4y11 + x6y8 + x8y5 + x10y2) << 272
        +   (x1y15 + x3y12 + x5y9 + x7y6 + x9y3) << 264
        +   (x2y13 + x4y10 + x6y7 + x8y4 + x10y1) << 256

        +   (x1y14 + x3y11 + x5y8 + x7y5 + x9y2) << 248
        +   (x0y15 + x2y12 + x4y9 + x6y6 + x8y3 + x10y0) << 240
        +   (x1y13 + x3y10 + x5y7 + x7y4 + x9y1) << 232
        +   (x2y11 + x0y14 + x4y8 + x6y5 + x8y2) << 224
        +   (x1y12 + x3y9 + x5y6 + x7y3 + x9y0) << 216
        +   (x0y13 + x2y10 + x4y7 + x6y4 + x8y1) << 208
        +   (x1y11 + x3y8 + x5y5 + x7y2) << 200
        +   (x0y12 + x2y9 + x4y6 + x6y3 + x8y0) << 192
        +   (x1y10 + x3y7 + x5y4 + x7y1) << 184
        +   (x0y11 + x2y8 + x4y5 + x6y2) << 176
        +   (x1y9 + x3y6 + x5y3 + x7y0) << 168
        +   (x0y10 + x2y7 + x4y4 + x6y1) << 160
        +   (x1y8 + x3y5 + x5y2) << 152
        +   (x0y9 + x2y6 + x4y3 + x6y0) << 144
        +   (x1y7 + x3y4 + x5y1) << 136
        +   (x0y8 + x2y5 + x4y2) << 128

        +   (x1y6 + x3y3 + x5y0) << 120
        +   (x0y7 + x2y4 + x4y1) << 112
        +   (x1y5 + x3y2) << 104
        +   (x0y6 + x2y3 + x4y0) << 96
        +   (x1y4 + x3y1) << 88
        +   (x2y2 + x0y5) << 80
        +   (x1y3 + x3y0) << 72
        +   (x0y4 + x2y1) << 64
        +   (x1y2) << 56
        +   (x0y3 + x2y0) << 48
        +   (x1y1) << 40
        +   (x0y2) << 32
        +   (x1y0) << 24
        +   (x0y1) << 16
        +   (x0y0)
    )
*/