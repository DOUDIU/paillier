module iddmm_top_tb();

parameter   K       =   256         ;// K bits in every group
parameter   N       =   16          ;// Number of groups
parameter   ADDR_W  =   $clog2(N)   ;

reg [K-1  :0]   wr_m1_                [0:3] = {
    256'h976ccf456fa1fb3bce136b8776f3a682ecd18b11b6a41b9bb3ef4fcae3ba221f,
    // 128'hecd18b11b6a41b9bb3ef4fcae3ba221f,
    128'hb885007f9c90c3f3beb79b92378fe7f,
    128'hb885007f9c90c3f3beb79b92378fe7f,
    128'hb885007f9c90c3f3beb79b92378fe7f
};

reg [K*N-1:0]   big_m                 [0:3] = {
    4096'hff5f4906fd176bc241535c78955d02f4d0acf376d736ae280077887200c758b7781b4432fa8baca2a81ad6fb0817051a00fccf8e15c63048681bcf8342b56433abd550affa489b289cd4f0482adce321c8cf4374ce15267692dfc8b0da108f4bb0e922d4a28402ef785c2516f6296486f8505ac3df05c0f953acce65e2dc5f1e59965ded73fa18ffb482ad1a2e5433d4df8211de12a3e7a71a1a084fed671fb11eeaf76f640c4fd549ea307b6622f798f027786e79232206de1507281d84c719209d408bc85f9ed2e1b82ecf72ff805a45221dc712c45a8dbc375e9b64227ec6b659a75fc5b5e051e776bcd9f4f6d82ebaff89a48c8494d6ed072372b846156af229994baab390ec57c00130255acc2cdf975783df4678153f0ca51b854425b1568b5b8b53239f50dd39fc53c3d41827a0687c435f6de5e98843def3fb7b0f7e701cdfb51517d6628392bd9291c16282556f5581766dd6a0a426a35312237399f93ad69502592c0f6d1864ba0b75600ee04cb406bcb833bc98527a0ac1249c6a918456b06f24611770c1708426b4d9041f7fe83be68fbc7018e461951d234ebf00227b4301911e24055c745203c888276f4db0c05f66514ae4e6b4bf4c8914e36c4a94bf57bf807dd40c7572d1a99c27d9f58af0877bb217c081d750d5edbe3c45eafc3ea6786560fa819873452cc8bffc7ab998ab70496b77fdadffb7ef2621,
    4096'h92d20837163355491353a40bfbed6afffb000939ca99e2dcb7e96c94d9e6ff1b54db47d62fa87283db4ef47e8119e2cb0d126f44ef110cd64d6493014fbee11fce25ad01515ed88bef11f595cc5b107aed44c3aecf42318a0e9dc2431934703c219abc2ee926037fbd46e2b2465b19b3110e3ccdbdfbe0daadefe22a725ef38bc2371fdc5e9cfb439ea6ac84b3e424e71cc3a263dc8cb4642042d01abe4e54416d821fae3e588950e16d5bdc76fc0629b4829eabad9ad1535fc322dc0ad791ca8a353157ab771cc0eafb621a07b0ce0998a65541754ffeedb756ff3ca3b606dea2b63fa2483a5dda07c17496f556f441e4c09fbb079cbbb8279c01fca24b56bf32e9902603d670439cee8a4f9730281ca7e736783300f69b64cce28fb565b99599758f8c8e5d58ce03af202cfe8d88092884f15b5a76578db8bf6a32cf7e2d78a758c60de9e6cf037bd2a6c7d22c670b8b384722fef18a9870588c1368f3c1f82caa709eff78cfdb2a3594bce3977875c0c30e464a5fc136225c7e206ba599b14ec856a9a230bca081331c969774eb112295c0670d4cb20723ceaa02e0ff4879a508052dad14c59f1787572686d68c51eb3ce8f505e141803ec18bc77c4986a7ea1dd24c13c7bb976496361ad38078e2daaf39f049a489793e2b46643b3eb3f168a3ad29eb4accb4ca422e7dd70e809f4ad5ed15d295f6765773bb5d851b3e81,
    4096'h92d20837163355491353a40bfbed6afffb000939ca99e2dcb7e96c94d9e6ff1b54db47d62fa87283db4ef47e8119e2cb0d126f44ef110cd64d6493014fbee11fce25ad01515ed88bef11f595cc5b107aed44c3aecf42318a0e9dc2431934703c219abc2ee926037fbd46e2b2465b19b3110e3ccdbdfbe0daadefe22a725ef38bc2371fdc5e9cfb439ea6ac84b3e424e71cc3a263dc8cb4642042d01abe4e54416d821fae3e588950e16d5bdc76fc0629b4829eabad9ad1535fc322dc0ad791ca8a353157ab771cc0eafb621a07b0ce0998a65541754ffeedb756ff3ca3b606dea2b63fa2483a5dda07c17496f556f441e4c09fbb079cbbb8279c01fca24b56bf32e9902603d670439cee8a4f9730281ca7e736783300f69b64cce28fb565b99599758f8c8e5d58ce03af202cfe8d88092884f15b5a76578db8bf6a32cf7e2d78a758c60de9e6cf037bd2a6c7d22c670b8b384722fef18a9870588c1368f3c1f82caa709eff78cfdb2a3594bce3977875c0c30e464a5fc136225c7e206ba599b14ec856a9a230bca081331c969774eb112295c0670d4cb20723ceaa02e0ff4879a508052dad14c59f1787572686d68c51eb3ce8f505e141803ec18bc77c4986a7ea1dd24c13c7bb976496361ad38078e2daaf39f049a489793e2b46643b3eb3f168a3ad29eb4accb4ca422e7dd70e809f4ad5ed15d295f6765773bb5d851b3e81,
    4096'h92d20837163355491353a40bfbed6afffb000939ca99e2dcb7e96c94d9e6ff1b54db47d62fa87283db4ef47e8119e2cb0d126f44ef110cd64d6493014fbee11fce25ad01515ed88bef11f595cc5b107aed44c3aecf42318a0e9dc2431934703c219abc2ee926037fbd46e2b2465b19b3110e3ccdbdfbe0daadefe22a725ef38bc2371fdc5e9cfb439ea6ac84b3e424e71cc3a263dc8cb4642042d01abe4e54416d821fae3e588950e16d5bdc76fc0629b4829eabad9ad1535fc322dc0ad791ca8a353157ab771cc0eafb621a07b0ce0998a65541754ffeedb756ff3ca3b606dea2b63fa2483a5dda07c17496f556f441e4c09fbb079cbbb8279c01fca24b56bf32e9902603d670439cee8a4f9730281ca7e736783300f69b64cce28fb565b99599758f8c8e5d58ce03af202cfe8d88092884f15b5a76578db8bf6a32cf7e2d78a758c60de9e6cf037bd2a6c7d22c670b8b384722fef18a9870588c1368f3c1f82caa709eff78cfdb2a3594bce3977875c0c30e464a5fc136225c7e206ba599b14ec856a9a230bca081331c969774eb112295c0670d4cb20723ceaa02e0ff4879a508052dad14c59f1787572686d68c51eb3ce8f505e141803ec18bc77c4986a7ea1dd24c13c7bb976496361ad38078e2daaf39f049a489793e2b46643b3eb3f168a3ad29eb4accb4ca422e7dd70e809f4ad5ed15d295f6765773bb5d851b3e81
};
reg [K*N-1:0]   big_x                 [0:3] = {
    4096'h7ffffffef380fcff68e38a9fcc30b4c64e94dbc4f2b03a88ae0650f51f46fe1f4f10ba102d77eb77c1547e0c40e6d7aeb05539c308ea01dafb6da33649210fab2cdd38a580091aaec64d74192431c00cce4f4c752498e88aaa5ccc010b2317db8e01cf660e1dc9ba01154024448965f8209721d391f8422ef2e1817ac4240be53bfc0f05b7336e172e271c9e9fcd38057746bbe8f5bb1907ab681ae012395e78e531f5291340108b4f8b182614a29fa0c7a44032229fe3fb3af01a5577cf335f318c1ecc70b613e7532ab85dc087c618020e949640cb14a3dbf634fa0b48f0098c9e9ee4861a5e6193f2a9241e28d1f4d3c9a8f11c460943dbd7b7b06f18fe75454e20593388dcaa8b98aabe293987d22e2725251d6ebf2729cde05db076ed775b7f369d1f9e1109812960b8b76e333bcca8aaa98931c2937cadb68a4ffc6c54eff9a6bcb77da76dc02fcb83167105319dd5a25f19d6ef0b214927120635e665afe46f681259247978d4a6853bb3cac03bc554d07003496f6b8b624bfec45f4cfb24acded0aeb074e8f70df1813ebb26bd5fe26be2a627684d793a8a052e3a9476a1d9697dd9e27beb4db7ad01eb8b0a3b5c7717d716ebd30727cc7786a17f09b04d6b94a56d9f70ac514e026f42834486e6a0852ce00808c7222cc02f90802ab22509fe316612d10d60359087ab7a23be6348b73f6704e6fde2ed070c500db0,4096'h7ffffffef380fcff68e38a9fcc30b4c64e94dbc4f2b03a88ae0650f51f46fe1f4f10ba102d77eb77c1547e0c40e6d7aeb05539c308ea01dafb6da33649210fab2cdd38a580091aaec64d74192431c00cce4f4c752498e88aaa5ccc010b2317db8e01cf660e1dc9ba01154024448965f8209721d391f8422ef2e1817ac4240be53bfc0f05b7336e172e271c9e9fcd38057746bbe8f5bb1907ab681ae012395e78e531f5291340108b4f8b182614a29fa0c7a44032229fe3fb3af01a5577cf335f318c1ecc70b613e7532ab85dc087c618020e949640cb14a3dbf634fa0b48f0098c9e9ee4861a5e6193f2a9241e28d1f4d3c9a8f11c460943dbd7b7b06f18fe75454e20593388dcaa8b98aabe293987d22e2725251d6ebf2729cde05db076ed775b7f369d1f9e1109812960b8b76e333bcca8aaa98931c2937cadb68a4ffc6c54eff9a6bcb77da76dc02fcb83167105319dd5a25f19d6ef0b214927120635e665afe46f681259247978d4a6853bb3cac03bc554d07003496f6b8b624bfec45f4cfb24acded0aeb074e8f70df1813ebb26bd5fe26be2a627684d793a8a052e3a9476a1d9697dd9e27beb4db7ad01eb8b0a3b5c7717d716ebd30727cc7786a17f09b04d6b94a56d9f70ac514e026f42834486e6a0852ce00808c7222cc02f90802ab22509fe316612d10d60359087ab7a23be6348b73f6704e6fde2ed070c500db0,4096'h6d2df7c8e9ccaab6ecac5bf40412950004fff6c635661d234816936b261900e4ab24b829d0578d7c24b10b817ee61d34f2ed90bb10eef329b29b6cfeb0411ee031da52feaea1277410ee0a6a33a4ef8512bb3c5130bdce75f1623dbce6cb8fc3de6543d116d9fc8042b91d4db9a4e64ceef1c33242041f2552101dd58da10c743dc8e023a16304bc6159537b4c1bdb18e33c5d9c23734b9bdfbd2fe541b1abbe927de051c1a776af1e92a4238903f9d64b7d615452652eaca03cdd23f5286e3575cacea85488e33f15049de5f84f31f66759aabe8ab0011248a900c35c49f9215d49c05db7c5a225f83e8b690aa90bbe1b3f6044f8634447d863fe035db4a940cd166fd9fc298fbc631175b068cfd7e35818c987ccff09649b331d704a9a466a668a707371a2a731fc50dfd3017277f6d77b0ea4a589a872474095cd3081d28758a739f2161930fc842d59382dd398f474c7b8dd010e75678fa773ec970c3e07d3558f6100873024d5ca6b431c68878a3f3cf1b9b5a03ec9dda381df945a664eb137a9565dcf435f7ecce369688b14eedd6a3f98f2b34df8dc3155fd1f00b7865af7fad252eb3a60e878a8d9792973ae14c3170afa1ebe7fc13e743883b6795815e22db3ec3844689b69c9e52c7f871d2550c60fb65b7686c1d4b99bc4c14c0e975c52d614b5334b35bdd18228f17f60b52a12ea2d6a0989a88c44a27ae4c17f,4096'h5b3c79741549edb3cfa435ec3658f9a1e3851eb89578184d3211d16d8301feac6e344ea52938af825d9c192e9cf7d8126f87a306462580c5f037719ee010123815dcbf70f2e7fd6c3ef5151072b1bdc841cf27ed8daed3f56798c4a3000e64ef02c6a96b4fe0ede0024b968f641550697364386ddb60e3d27074c78f32d3f50b7df51c860725c40420aed07295ccb45d5c2b508e6f5c56d0502b1cd8078342da541b93752507d20f04315e90d19875541808eb9dbc3278b8ed2d0d4c28891db296a74f3b76fd8b81a7cedc4f439efa159ed76724cc551be0d1f05d0f35739d5f23ba6b560ea8567457fb669ca9eef8550ebeaace53ce1c866ae4e6de6b6a4d617bb77ca72fda2cbe4bddae2a0983a133dd3af895b747de0d5efbadb2e97da51e8d4a1746321a4e7380551a8b40d0c80aa9b8e2aa281e2fae18b783b584fd2efd52d3a208a3bea1da7a0750317f3e12d67646849cb97ae5508cabe2bfacaaaba01372d38f22744b67055900556784824f329626655d0b7792d8ab80c08a0f0e33c7df6b52709117e4ffbcf65492de2691d1271c8c29e2d3d845f6a8c43cccca8ef05c2aff8ecc15e52e32151090d9d6b63b437a88e9ab12a1a42f5a0639d66552b80c89333a8c2ae1ad7bd9d40bcbbb7445954b4615d636e323e7c7d8d1b19d16320069e41ca37f938b1a4b17e837cd05e5c4cab9ed9db2e5649e0dddb42fdf91
};
reg [K*N-1:0]   big_y                 [0:3] = {
    4096'h9ffff4f73caff09ff67fc82fe8f5988fe76cff5b4241f1f3f3f4ccb35f29fff573f617bc077c80165ec5270c0b863fc231ae96dd5d933e9a98abdaf3d6e852e98149945ab1a9a90e38e07c3017c1273b18598d87b59a289de9d7c5bc5c6f64cccdbcbec42c289c8b1b799f8454cba6b89e5976a84c19217d64ddde5af42e37ab465928d068deaa3a0270b8d062dbe0b737667c3afd065871532081e72bc1f79e1d7ebd1fb933ec3555a8e986f949f72ca11bc2fbe4c704b20838c68b707d9f3db1d8ae45b44b6bd36a58bfbf7d565347a6c6e20130c84f1bad77f6251e81dfb6ffa9a508d64db7d2fe48b5e4ebe68e7c8d62cdf5ab1c2ca8c2d2e835a1423acbef65956c980dfb62b3a405b9efbc93283d5071c2129b831481c537cc5be8f1d2723f1168f797bde736c1f73054d7d0dc97538fba25bb3e38703934d8fc46ad22eb23ea409184c3dba8241efc92ce5a6728f4385da637bc23ef7acb506d0543804ae7d660926a82406f9d3206376d5454466ecde2246a125c99aebdf16743d55cfb1c4ab0fdb8387320d541a94e3c5aa6038466eaa18682a163d571db3214de448b3d4d7a632bc60f0a524a041cd6e72a75dbc9f6bb63743df3c3c0d4649a28bd0bbeee569182303a66b830a2273b8df05c712adadf2bcb75244a66826265da778e0c3b45a20d6c962fd203e708ff62dd29b9edd90f2afd2bfe92014968e4396a,4096'h915f94ab9c50ca4ab4eeed592a9beaa5ad6f3ab8cde33356263b7ca1cd6327f93abe0f5f621642eb55318e74137d0b258ebc8b10a00cab3ffe67b8e78a16a98e4ddb4c9ac0c0a08302a84f682ca131a477edce6c0888a7d3b0aa71c00185447b162a3b903f9853566121da8222821f4429e054b3919b6c6c038207f135accb78acd282aca5f291fca5ea2cc846ae54dffe7b604b0be2fe402bcb234c62e040177915fd96957f012fc6c3c43fa5b2e41107252f907ab98a98c4d0dd09e90ef2e0f4a75b8a7d8b166e180cb21a76528f23f9a7752b5ac26ac1e8c15c514343b84b3b1450e77af95bdf8148328d73d65a6cd4479f00aaf1fe6a7641a67c0515e8f6e169cc22bf64c781c30d0a498b07001a95d7776b9beb874091aeaabc1594693fd8ea828ac8251e7835669e4adb373a0f24428720ad662853fbb3f3f4d95cf52de704570cefbc67502abb2837ea155c3df5e87eb6400b55d7ec696534b23ed3774ed73d9fc2788919bf9d984c670019bd4d0a8c0ba1be9c46ce46811a7f8fbaea6e74eb0c8d4989c5f7f7ba424a380576979df18527249a66e10251090d2bad6a25fa45d9a2ce695e98e2ae4f3b06c5f3c72909e099111c79ca5511174ff3fb35f3e16d1d8e50675156b0f608a0c7d82b62d7b109a4be8fceb700f50b47c35664ce312818a6f6c0b2ff78a1ac2de5674a4fcaa08ceba5ea9d842695dd79db7aa0,
    4096'h6d2df7c8e9ccaab6ecac5bf40412950004fff6c635661d234816936b261900e4ab24b829d0578d7c24b10b817ee61d34f2ed90bb10eef329b29b6cfeb0411ee031da52feaea1277410ee0a6a33a4ef8512bb3c5130bdce75f1623dbce6cb8fc3de6543d116d9fc8042b91d4db9a4e64ceef1c33242041f2552101dd58da10c743dc8e023a16304bc6159537b4c1bdb18e33c5d9c23734b9bdfbd2fe541b1abbe927de051c1a776af1e92a4238903f9d64b7d615452652eaca03cdd23f5286e3575cacea85488e33f15049de5f84f31f66759aabe8ab0011248a900c35c49f9215d49c05db7c5a225f83e8b690aa90bbe1b3f6044f8634447d863fe035db4a940cd166fd9fc298fbc631175b068cfd7e35818c987ccff09649b331d704a9a466a668a707371a2a731fc50dfd3017277f6d77b0ea4a589a872474095cd3081d28758a739f2161930fc842d59382dd398f474c7b8dd010e75678fa773ec970c3e07d3558f6100873024d5ca6b431c68878a3f3cf1b9b5a03ec9dda381df945a664eb137a9565dcf435f7ecce369688b14eedd6a3f98f2b34df8dc3155fd1f00b7865af7fad252eb3a60e878a8d9792973ae14c3170afa1ebe7fc13e743883b6795815e22db3ec3844689b69c9e52c7f871d2550c60fb65b7686c1d4b99bc4c14c0e975c52d614b5334b35bdd18228f17f60b52a12ea2d6a0989a88c44a27ae4c17f,
    4096'h5b3c79741549edb3cfa435ec3658f9a1e3851eb89578184d3211d16d8301feac6e344ea52938af825d9c192e9cf7d8126f87a306462580c5f037719ee010123815dcbf70f2e7fd6c3ef5151072b1bdc841cf27ed8daed3f56798c4a3000e64ef02c6a96b4fe0ede0024b968f641550697364386ddb60e3d27074c78f32d3f50b7df51c860725c40420aed07295ccb45d5c2b508e6f5c56d0502b1cd8078342da541b93752507d20f04315e90d19875541808eb9dbc3278b8ed2d0d4c28891db296a74f3b76fd8b81a7cedc4f439efa159ed76724cc551be0d1f05d0f35739d5f23ba6b560ea8567457fb669ca9eef8550ebeaace53ce1c866ae4e6de6b6a4d617bb77ca72fda2cbe4bddae2a0983a133dd3af895b747de0d5efbadb2e97da51e8d4a1746321a4e7380551a8b40d0c80aa9b8e2aa281e2fae18b783b584fd2efd52d3a208a3bea1da7a0750317f3e12d67646849cb97ae5508cabe2bfacaaaba01372d38f22744b67055900556784824f329626655d0b7792d8ab80c08a0f0e33c7df6b52709117e4ffbcf65492de2691d1271c8c29e2d3d845f6a8c43cccca8ef05c2aff8ecc15e52e32151090d9d6b63b437a88e9ab12a1a42f5a0639d66552b80c89333a8c2ae1ad7bd9d40bcbbb7445954b4615d636e323e7c7d8d1b19d16320069e41ca37f938b1a4b17e837cd05e5c4cab9ed9db2e5649e0dddb42fdf91
};
reg [K*N-1:0]   iddmm_result_confirm  [0:3] = {
    4096'h47a205a79ebd89394649f7942601cf1ea095b448c7c5054237b6657725c08e56a4edc79ccc6c9f83c801b2098246b1f3eb991a4634cd993b221dbd3b9b0fecacf4ffd56189592bd5c668399022496765705a0c9dcfb5da9d79c0e001f14ef78f2c895ab0bbf9b5ea5021fc316a0aa7b17b4b2c8ef8723f2ac3698ec872875b69ceaa84e184c4481bfa53cb2d99f029439fe9564393756f591dd20c30984eddbeb44e9e5104dbc64fbf4bc88319115cf49b21eb137f5a1576ea5819224800f2977285a611de039cd1049a62cb3f4e67d9c65dc48af76555819e57712018989b6f46fd06e477938b79ee8246fd27349abef24f5738173925dbfbace3f264e7edec8cb836900e60b5a59af3c56f14d8953d3411f9bad910846eff8d9f1796723722a88dda362be3abfec27f67cc32bdc7d41e2848d56d9d91cd754765a3e5a171e5964d862cc64a3437e1a35a997fe47ead24c2e5823ef70acc9ac946f3f00bc0177146d68369a8b607a72392b9dea6ee7477baaaa4a50106aa648ff4f4da63d8f3306116466a289c0d9927606cd104cfe8e3ae65849bbe124fc61ebf289c2f5cf1399aa5bf08aeef91fb4b542ce253a87b89ec9ce0a4be3914a67d44b6a8fa5678d8e8d1185ab86cac8472aad50c039115b61790a2c7dbe2e7bdc94990f1d6bb0aa0a5613d7387216fe18c1a0fe6b9388bf708ee9a9074da10a576774987b41f6a,
    4096'h23e5cecd1b969f69f024855e671bb4d40fad9200b83f289b72f43a28c4e12884c14f8754d535d4ed623f2689fd2b3b7905874e6cfb0d03baf027b9ccb1cce4cee606a091db56ed2dfa876528a5feef5e0839b6082a5e261eef12ce67dd4b0fafb6627ae7cc0c339e5b77f52d2b2be2d10ad3470e9a3dd062e8a7e2c62eaaf3703071434f77002c5020c0f1bc025858f26c808182366c83afc05e9bc6e2d8d6b98dd559eb2c91414169d545ac449404e3e7fdfe3716add38bb1defbc9d6ed663c266a34562aa9dc34ad0dd319391e6ae7ce1a2882f72d8b41860e95e08a78e290e9ef30f43438d836ec229d4d6e33478901498f51535f4bbdb8e2b4e1c59e38decb8424416840b8da4a12d5704a2ece92425151ae37e45edc677aa7402d50ee3284c4e1c9fdc1a826a2eb241a9a95553af156511f4c1639422c134c49ee0091e2799bac77e6bf069a2cefae4a251ed0d49256285c3540ad6194bfe68d4dc3e5d47a537228a9f214d60b18308c8ca1194bec2c500daec1abaefb528f18dccb96420c1b020a488553b8807baa6e16d72c61cf8fb63b3665317441036d3c0ee61924a742adee2cb0678d93244f79d6cb566ae7977e425d6ae5853fc062f9890f7c67a00db107cd3f0c98cf97a0f7efa95d9e8fe00afbf5b0cae721055edd7ab577bdb6c5a0ffa814a24fd759556fb81f23c036d1c31cfca5a1d6c1e0c2d56ed98f27,
    4096'h6d2df7c8e9ccaab6ecac5bf40412950004fff6c635661d234816936b261900e4ab24b829d0578d7c24b10b817ee61d34f2ed90bb10eef329b29b6cfeb0411ee031da52feaea1277410ee0a6a33a4ef8512bb3c5130bdce75f1623dbce6cb8fc3de6543d116d9fc8042b91d4db9a4e64ceef1c33242041f2552101dd58da10c743dc8e023a16304bc6159537b4c1bdb18e33c5d9c23734b9bdfbd2fe541b1abbe927de051c1a776af1e92a4238903f9d64b7d615452652eaca03cdd23f5286e3575cacea85488e33f15049de5f84f31f66759aabe8ab0011248a900c35c49f9215d49c05db7c5a225f83e8b690aa90bbe1b3f6044f8634447d863fe035db4a940cd166fd9fc298fbc631175b068cfd7e35818c987ccff09649b331d704a9a466a668a707371a2a731fc50dfd3017277f6d77b0ea4a589a872474095cd3081d28758a739f2161930fc842d59382dd398f474c7b8dd010e75678fa773ec970c3e07d3558f6100873024d5ca6b431c68878a3f3cf1b9b5a03ec9dda381df945a664eb137a9565dcf435f7ecce369688b14eedd6a3f98f2b34df8dc3155fd1f00b7865af7fad252eb3a60e878a8d9792973ae14c3170afa1ebe7fc13e743883b6795815e22db3ec3844689b69c9e52c7f871d2550c60fb65b7686c1d4b99bc4c14c0e975c52d614b5334b35bdd18228f17f60b52a12ea2d6a0989a88c44a27ae4c17f,
    4096'h103588031a2919264e97c60a2aad4c1d5efda770b830222207b2f9743a8e3aee4ccb4213ff81f16c6fe41363ff4256fa808ff2359fbaaefa5dc7e12c9198058e6912ebc92add92cef48fd1b2310c03419f206faedbee0b78b598f82eae3209286bf91852db03228a26a94f04400a3236b46503b792c73258b3f290871e138ef22ee4e3eb365e60674d51674d3ef3218312c02400e6348831aa54694506222be49eb73a2d09e428ba97c04d5c12bf9be526706a8dd7071ab74a7a283309f19ec9c87c63cd6e0f95c909243cbbf56fb20e96e5cf30d863f94e574eb5ac6bef6d2e8d95054d64f34e31570256eeeb092f2c23dc9be8794fbf29af45bf9bc732941385e88b1ca6d2a506ce8826387435d097d60e2f152f673f19c26a22f18fe95e7535339860202130531cd4d84272963b9f9521eb5f30f9dd74e17e80d2963c0a6712a0302ce3d78cae15d162513175bb129a22ab7a33db808f24dd4fcbb426f10dbc4a1a90ad9a11a70a0acf9cda7d099ef88338672d41e66fc63f44f3fc770858e802939fc6b8888ad8a276b92d7bf79d7f1a7e519caa5060a84d1e86c1dac2d76bb5f387fa1ec81b0587b37bb5d2d35ac83437c8be7edd4fa6934874f1d9164832c6bb2c6c7a804fc1996d86ffbaf5b8fb29607dc0d875feb37cc7990d5b1a75488de47453202db9c7dfc669589399598806cca2db96e82ea458f2f4bb040b96
};

reg [K*N-1:0]   iddmm_result = 0; 

reg clk = 0;
reg rst_n = 0;
always #5 clk = ~clk;
initial #30 rst_n = 1;


reg     [2          :0]     wr_ena          ;
reg     [ADDR_W-1   :0]     wr_addr         ;
reg     [K-1        :0]     wr_x            ;
reg     [K-1        :0]     wr_y            ;
reg     [K-1        :0]     wr_m            ;
reg     [K-1        :0]     wr_m1           ;

reg                         task_req        ;
wire                        task_end        ;
wire                        task_grant      ;
wire    [K-1        :0]     task_res        ;

task single_request(input num);
    integer i;

    for(i = 0; i < N; i = i + 1) begin
        wr_ena      <=  3'b111;
        wr_addr     <=  i;
        wr_x        <=  big_x [num][i*K +: K];
        wr_y        <=  big_y [num][i*K +: K];
        wr_m        <=  big_m [num][i*K +: K];
        wr_m1       <=  wr_m1_[num];
        @(posedge clk);
    end

    @(posedge clk);
    task_req    <=  1;
    @(posedge clk);
    task_req    <=  0;

    wait(task_grant);
    for(i = 0; i < N; i = i + 1) begin
        @(posedge clk);
        iddmm_result[i*K +: K]   <=  task_res;
    end
    @(posedge clk);
    assert(iddmm_result ==  iddmm_result_confirm[num])
        $display("result is correct!");
    else begin
        $display("result is wrong!");
        $display("iddmm_result = %h", iddmm_result); 
        $display("iddmm_result_confirm = %h", iddmm_result_confirm[num]); 
    end
endtask


initial begin
    wr_ena      <=  0;
    wr_addr     <=  0;
    wr_x        <=  0;
    wr_y        <=  0;
    wr_m        <=  0;
    wr_m1       <=  0;
    task_req    <=  0;
    @(posedge rst_n);
    for(int i = 0; i < 1; i = i + 1) begin
        single_request(i);
    end
    $stop;
end

iddmm_top #(
        .K              (K          )
    ,   .N              (N          )
)iddmm_top_inst(
        .clk            (clk        )
    ,   .rst_n          (rst_n      )

    ,   .wr_ena         (wr_ena     )
    ,   .wr_addr        (wr_addr    )
    ,   .wr_x           (wr_x       )
    ,   .wr_y           (wr_y       )
    ,   .wr_m           (wr_m       )
    ,   .wr_m1          (wr_m1      )

    ,   .task_req       (task_req   )
    ,   .task_end       (task_end   )
    ,   .task_grant     (task_grant )
    ,   .task_res       (task_res   )
);


endmodule