module L_func_top #(
        parameter K       = 128
    ,   parameter N       = 32
)(
        input               clk
    ,   input               rst_n

    ,   input               task_start

    ,   input   [K-1:0]     L_x
    ,   input               L_x_valid

    ,   output  [K-1:0]     L_out
    ,   output              L_out_valid
);

























































endmodule